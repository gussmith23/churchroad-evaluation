module mul_0_stage_unsigned_16_16_16_bit(input [15:0] a, b, output [15:0] out);
  assign out = a * b;
endmodule